library verilog;
use verilog.vl_types.all;
entity LZE_vlg_check_tst is
    port(
        result          : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end LZE_vlg_check_tst;
