library verilog;
use verilog.vl_types.all;
entity RED_vlg_vec_tst is
end RED_vlg_vec_tst;
