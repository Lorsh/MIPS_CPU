library verilog;
use verilog.vl_types.all;
entity RED is
    port(
        input1          : in     vl_logic_vector(31 downto 0);
        result          : out    vl_logic_vector(7 downto 0)
    );
end RED;
