library verilog;
use verilog.vl_types.all;
entity UZE_vlg_vec_tst is
end UZE_vlg_vec_tst;
