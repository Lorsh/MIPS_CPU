library verilog;
use verilog.vl_types.all;
entity LZE_vlg_vec_tst is
end LZE_vlg_vec_tst;
