LIBRARY ieee; 
USE ieee.std_logic_1164.ALL;  
USE ieee.std_logic_arith.ALL;  
USE ieee.std_logic_unsigned.ALL; 

ENTITY mux_8to1 IS 
PORT(
in0,in1,in2,in3,in4,in5,in6,in7		:IN STD_LOGIC_VECTOR(31 DOWNTO 0);  
selector     : IN STD_LOGIC_VECTOR( 2 DOWNTO 0);  
result   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));  
END mux_8to1; 


ARCHITECTURE description OF mux_8to1 IS
BEGIN
	process (in0,in1,in2,in3,in4,in5,in6,in7) 
		BEGIN
			case selector is
				when "000" =>
					result <= in0;
				when 	"001" =>
					result <= in1;
				when "010" =>
					result <= in2;
				when "011" =>
					result <= in3;
				when 	"100" =>
					result <= in4;
				when "101" =>
					result <= in5;
				when "110" =>
					result <= in6;
				when 	"111" =>
					result <= in7;
				when others => result <= "ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ"; --in case some weird input comes in that is not one of the above
				
			end case;
		end process;
END description;